-- Scrolls the game state and generates new notes to play

--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.numeric_std.all;
--use IEEE.std_logic_unsigned.all;

-- This should do something to generate a new 1 or 0 on top of the string. Needs to be random?